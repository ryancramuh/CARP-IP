`ifndef CLK_PARAMS_SVH
`define CLK_PARAMS_SVH

parameter CLKS_PER_BIT_100MHZ 868
parameter CLKS_PER_BIT_10MHZ 87

`endif
